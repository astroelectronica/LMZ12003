.title KiCad schematic
.include "C:/AE/LMZ12003/_models/C2012X7R2A223K125AE_p.mod"
.include "C:/AE/LMZ12003/_models/C3216X5R0J107M160AB_p.mod"
.include "C:/AE/LMZ12003/_models/C3216X7R1H105K160AE_p.mod"
.include "C:/AE/LMZ12003/_models/C3225X5R1H106K250AB_p.mod"
.include "C:/AE/LMZ12003/_models/LMZ12003_TRANS.LIB"
XU7 VDD 0 C3216X5R0J107M160AB_p
XU3 VDD /FB C2012X7R2A223K125AE_p
R4 VDD /FB {RFBT}
R6 VDD 0 {RLOAD}
XU5 VDD 0 C3216X7R1H105K160AE_p
R2 /EN 0 {RENB}
R1 VCC /EN {RENT}
XU1 VCC /RON /EN 0 /SS /FB VDD LMZ12003_TRANS
R3 /RON VCC {RON}
XU4 VCC 0 C3216X7R1H105K160AE_p
XU6 VCC 0 C3225X5R1H106K250AB_p
XU2 /SS 0 C2012X7R2A223K125AE_p
R5 /FB 0 {RFBB}
V1 VCC 0 {VIN}
.end
